module char_gen (
    input [5:0] char, 
    input [2:0] row,
    output reg [7:0] pixels
);

/* 
    ENCODING    CHARACTER
           0            0
           1            1
           2            2
           3            3
           4            4
           5            5
           6            6
           7            7
           8            8
           9            9
          10            A
          11            B
          12            C
          13            D
          14            E
          15            F
          16            G
          17            H
          18            I
          19            J
          20            K
          21            L
          22            M  
          23            N
          24            O
          25            P
          26            Q
          27            R
          28            S
          29            T
          30            U
          31            V
          32            W
          33            X
          34            Y
          35            Z
          36            !
          37            ?
          38           ' ' (space)
*/

always @(*) begin 
    case ({char,row})
        10'b000000_000: pixels = 8'b01111100; //  XXXXX  |
        10'b000000_001: pixels = 8'b11000110; // XX   XX |
        10'b000000_010: pixels = 8'b11000110; // XX   XX |
        10'b000000_011: pixels = 8'b11000110; // XX   XX |
        10'b000000_100: pixels = 8'b11000110; // XX   XX |
        10'b000000_101: pixels = 8'b11000110; // XX   XX |
        10'b000000_110: pixels = 8'b01111100; //  XXXXX  |
        10'b000000_111: pixels = 8'b00000000; // ________|

        10'b000001_000: pixels = 8'b00011000; //    XX   |
        10'b000001_001: pixels = 8'b00111000; //   XXX   |
        10'b000001_010: pixels = 8'b00011000; //    XX   |
        10'b000001_011: pixels = 8'b00011000; //    XX   |
        10'b000001_100: pixels = 8'b00011000; //    XX   |
        10'b000001_101: pixels = 8'b00011000; //    XX   |
        10'b000001_110: pixels = 8'b00111110; //  XXXXXX |
        10'b000001_111: pixels = 8'b00000000; // ________|

        10'b000010_000: pixels = 8'b01111100; //  XXXXX  |
        10'b000010_001: pixels = 8'b11101110; // XXX XXX |
        10'b000010_010: pixels = 8'b00001110; //     XXX |
        10'b000010_011: pixels = 8'b00011100; //    XXX  |
        10'b000010_100: pixels = 8'b00111000; //   XXX   |
        10'b000010_101: pixels = 8'b01110000; //  XXX    |
        10'b000010_110: pixels = 8'b11111110; // XXXXXXX |
        10'b000010_111: pixels = 8'b00000000; // ________|

        10'b000011_000: pixels = 8'b01111100; //  XXXXX  |
        10'b000011_001: pixels = 8'b11000110; // XX   XX |
        10'b000011_010: pixels = 8'b00000110; //      XX |
        10'b000011_011: pixels = 8'b00011100; //    XXX  |
        10'b000011_100: pixels = 8'b00000110; //      XX |
        10'b000011_101: pixels = 8'b11000110; // XX   XX |
        10'b000011_110: pixels = 8'b01111100; //  XXXXX  |
        10'b000011_111: pixels = 8'b00000000; // ________|

        10'b000100_000: pixels = 8'b01100110; //  XX  XX |
        10'b000100_001: pixels = 8'b01100110; //  XX  XX |
        10'b000100_010: pixels = 8'b01100110; //  XX  XX |
        10'b000100_011: pixels = 8'b01111110; //  XXXXXX |
        10'b000100_100: pixels = 8'b00000110; //      XX |
        10'b000100_101: pixels = 8'b00000110; //      XX |
        10'b000100_110: pixels = 8'b00000110; //      XX |
        10'b000100_111: pixels = 8'b00000000; // ________|

        10'b000101_000: pixels = 8'b11111110; // XXXXXXX |
        10'b000101_001: pixels = 8'b11000000; // XX      |
        10'b000101_010: pixels = 8'b11111000; // XXXXX   |
        10'b000101_011: pixels = 8'b00000110; //      XX |
        10'b000101_100: pixels = 8'b00000110; //      XX |
        10'b000101_101: pixels = 8'b11001100; // XX  XX  |
        10'b000101_110: pixels = 8'b11111000; // XXXXX   |
        10'b000101_111: pixels = 8'b00000000; // ________|

        10'b000110_000: pixels = 8'b11111110; // XXXXXXX |
        10'b000110_001: pixels = 8'b11000000; // XX      |
        10'b000110_010: pixels = 8'b11000000; // XX      |
        10'b000110_011: pixels = 8'b11111110; // XXXXXXX |
        10'b000110_100: pixels = 8'b11000110; // XX   XX |
        10'b000110_101: pixels = 8'b11000110; // XX   XX |
        10'b000110_110: pixels = 8'b11111110; // XXXXXXX |
        10'b000110_111: pixels = 8'b00000000; // ________|

        10'b000111_000: pixels = 8'b11111100; // XXXXXX  |
        10'b000111_001: pixels = 8'b11000110; // XX  XX  |
        10'b000111_010: pixels = 8'b00000110; //     XX  |
        10'b000111_011: pixels = 8'b00001100; //    XX   |
        10'b000111_100: pixels = 8'b00011000; //   XX    |
        10'b000111_101: pixels = 8'b00011000; //   XX    |
        10'b000111_110: pixels = 8'b00011000; //   XX    |
        10'b000111_111: pixels = 8'b00000000; // ________|

        10'b001000_000: pixels = 8'b01111100; //  XXXXX  |
        10'b001000_001: pixels = 8'b11000110; // XX   XX |
        10'b001000_010: pixels = 8'b11000110; // XX   XX |
        10'b001000_011: pixels = 8'b01111100; //  XXXXX  |
        10'b001000_100: pixels = 8'b11000110; // XX   XX |
        10'b001000_101: pixels = 8'b11000110; // XX   XX |
        10'b001000_110: pixels = 8'b01111100; //  XXXXX  |
        10'b001000_111: pixels = 8'b00000000; // ________|

        10'b001001_000: pixels = 8'b01111100; //  XXXXX  |
        10'b001001_001: pixels = 8'b11000110; // XX   XX |
        10'b001001_010: pixels = 8'b11000110; // XX   XX |
        10'b001001_011: pixels = 8'b01111110; //  XXXXXX |
        10'b001001_100: pixels = 8'b00000110; //      XX |
        10'b001001_101: pixels = 8'b00001100; //     XX  |
        10'b001001_110: pixels = 8'b00011000; //    XX   |
        10'b001001_111: pixels = 8'b00000000; // ________|

        10'b001010_000: pixels = 8'b00111000; //   XXX   |
        10'b001010_001: pixels = 8'b01101100; //  XX XX  |
        10'b001010_010: pixels = 8'b11000110; // XX   XX |
        10'b001010_011: pixels = 8'b11000110; // XX   XX |
        10'b001010_100: pixels = 8'b11111110; // XXXXXXX |
        10'b001010_101: pixels = 8'b11000110; // XX   XX |
        10'b001010_110: pixels = 8'b11000110; // XX   XX |
        10'b001010_111: pixels = 8'b00000000; // ________|

        
